
module Instr_Mem(A,rst,RD );
input [31:0] A;
input rst;
output [31:0]RD;

reg [31:0]Mem [1023:0];

assign RD=(rst==1'b0)?32'h00000000:Mem[A[31:2]];
initial begin
//Mem[0]=32'hFFC4A303;
//Mem[1]=32'h00832383;
Mem[0]=32'h00500293;
Mem[1]=32'h00300313;

Mem[2]=32'h006283B3;
Mem[3]=32'h00002403;
Mem[4]=32'h00100493;
Mem[5]=32'h00940533;
end 
/*initial begin
$readmemh("memfile.hex",Mem);
end*/
endmodule
